library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;

    use work.Types.all;

entity FirstRom is
    port (
        clk: in  std_logic;
        addressX: in integer range 0 to 27; 
        addressY: in integer range 0 to 27;
        addressZ: in integer range 0 to 2;

        output: out unsigned(15 downto 0)
    );
end entity;

architecture rtl of FirstRom is

begin
    process(all)
    begin
        if rising_edge(clk) then 
            case addressX is
                when 0 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 1 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 2 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 3 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 4 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 5 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 6 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 7 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 8 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 9 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000100001101";
                                when 1 =>
                                    output <= "0000000100001101";
                                when others =>
                                    output <= "0000000100001101";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000010110100";
                                when 1 =>
                                    output <= "0000000010110100";
                                when others =>
                                    output <= "0000000010110100";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 10 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000010000";
                                when 1 =>
                                    output <= "0000000000010000";
                                when others =>
                                    output <= "0000000000010000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000101100001";
                                when 1 =>
                                    output <= "0000000101100001";
                                when others =>
                                    output <= "0000000101100001";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001011011110";
                                when 1 =>
                                    output <= "0000001011011110";
                                when others =>
                                    output <= "0000001011011110";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111111011";
                                when 1 =>
                                    output <= "0000001111111011";
                                when others =>
                                    output <= "0000001111111011";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111111011";
                                when 1 =>
                                    output <= "0000001111111011";
                                when others =>
                                    output <= "0000001111111011";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111011011";
                                when 1 =>
                                    output <= "0000001111011011";
                                when others =>
                                    output <= "0000001111011011";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000101111001";
                                when 1 =>
                                    output <= "0000000101111001";
                                when others =>
                                    output <= "0000000101111001";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000100000";
                                when 1 =>
                                    output <= "0000000000100000";
                                when others =>
                                    output <= "0000000000100000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110100101";
                                when 1 =>
                                    output <= "0000000110100101";
                                when others =>
                                    output <= "0000000110100101";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101011011";
                                when 1 =>
                                    output <= "0000001101011011";
                                when others =>
                                    output <= "0000001101011011";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110100011";
                                when 1 =>
                                    output <= "0000001110100011";
                                when others =>
                                    output <= "0000001110100011";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 11 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001001000";
                                when 1 =>
                                    output <= "0000000001001000";
                                when others =>
                                    output <= "0000000001001000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101011111";
                                when 1 =>
                                    output <= "0000001101011111";
                                when others =>
                                    output <= "0000001101011111";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101011011";
                                when 1 =>
                                    output <= "0000001101011011";
                                when others =>
                                    output <= "0000001101011011";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000111110001";
                                when 1 =>
                                    output <= "0000000111110001";
                                when others =>
                                    output <= "0000000111110001";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000010110100";
                                when 1 =>
                                    output <= "0000000010110100";
                                when others =>
                                    output <= "0000000010110100";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101011011";
                                when 1 =>
                                    output <= "0000001101011011";
                                when others =>
                                    output <= "0000001101011011";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001100000111";
                                when 1 =>
                                    output <= "0000001100000111";
                                when others =>
                                    output <= "0000001100000111";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000011010000";
                                when 1 =>
                                    output <= "0000000011010000";
                                when others =>
                                    output <= "0000000011010000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001100111011";
                                when 1 =>
                                    output <= "0000001100111011";
                                when others =>
                                    output <= "0000001100111011";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001100111111";
                                when 1 =>
                                    output <= "0000001100111111";
                                when others =>
                                    output <= "0000001100111111";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110101001";
                                when 1 =>
                                    output <= "0000000110101001";
                                when others =>
                                    output <= "0000000110101001";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 12 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000011000";
                                when 1 =>
                                    output <= "0000000000011000";
                                when others =>
                                    output <= "0000000000011000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110011101";
                                when 1 =>
                                    output <= "0000000110011101";
                                when others =>
                                    output <= "0000000110011101";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110101011";
                                when 1 =>
                                    output <= "0000001110101011";
                                when others =>
                                    output <= "0000001110101011";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101010011";
                                when 1 =>
                                    output <= "0000001101010011";
                                when others =>
                                    output <= "0000001101010011";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000011111100";
                                when 1 =>
                                    output <= "0000000011111100";
                                when others =>
                                    output <= "0000000011111100";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000010100";
                                when 1 =>
                                    output <= "0000000000010100";
                                when others =>
                                    output <= "0000000000010100";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110001111";
                                when 1 =>
                                    output <= "0000001110001111";
                                when others =>
                                    output <= "0000001110001111";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001010011110";
                                when 1 =>
                                    output <= "0000001010011110";
                                when others =>
                                    output <= "0000001010011110";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000100";
                                when 1 =>
                                    output <= "0000000000000100";
                                when others =>
                                    output <= "0000000000000100";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000100000001";
                                when 1 =>
                                    output <= "0000000100000001";
                                when others =>
                                    output <= "0000000100000001";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110011011";
                                when 1 =>
                                    output <= "0000001110011011";
                                when others =>
                                    output <= "0000001110011011";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111101011";
                                when 1 =>
                                    output <= "0000001111101011";
                                when others =>
                                    output <= "0000001111101011";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101111111";
                                when 1 =>
                                    output <= "0000001101111111";
                                when others =>
                                    output <= "0000001101111111";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000010110100";
                                when 1 =>
                                    output <= "0000000010110100";
                                when others =>
                                    output <= "0000000010110100";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000010000";
                                when 1 =>
                                    output <= "0000000000010000";
                                when others =>
                                    output <= "0000000000010000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 13 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000111100101";
                                when 1 =>
                                    output <= "0000000111100101";
                                when others =>
                                    output <= "0000000111100101";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001010100110";
                                when 1 =>
                                    output <= "0000001010100110";
                                when others =>
                                    output <= "0000001010100110";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001001000";
                                when 1 =>
                                    output <= "0000000001001000";
                                when others =>
                                    output <= "0000000001001000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000100011101";
                                when 1 =>
                                    output <= "0000000100011101";
                                when others =>
                                    output <= "0000000100011101";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111100011";
                                when 1 =>
                                    output <= "0000001111100011";
                                when others =>
                                    output <= "0000001111100011";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000100111001";
                                when 1 =>
                                    output <= "0000000100111001";
                                when others =>
                                    output <= "0000000100111001";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001001000110";
                                when 1 =>
                                    output <= "0000001001000110";
                                when others =>
                                    output <= "0000001001000110";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110001111";
                                when 1 =>
                                    output <= "0000001110001111";
                                when others =>
                                    output <= "0000001110001111";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110100001";
                                when 1 =>
                                    output <= "0000000110100001";
                                when others =>
                                    output <= "0000000110100001";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000101100";
                                when 1 =>
                                    output <= "0000000000101100";
                                when others =>
                                    output <= "0000000000101100";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 14 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110001001";
                                when 1 =>
                                    output <= "0000000110001001";
                                when others =>
                                    output <= "0000000110001001";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111011111";
                                when 1 =>
                                    output <= "0000001111011111";
                                when others =>
                                    output <= "0000001111011111";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110110101";
                                when 1 =>
                                    output <= "0000000110110101";
                                when others =>
                                    output <= "0000000110110101";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000010000";
                                when 1 =>
                                    output <= "0000000000010000";
                                when others =>
                                    output <= "0000000000010000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000111000";
                                when 1 =>
                                    output <= "0000000000111000";
                                when others =>
                                    output <= "0000000000111000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110000011";
                                when 1 =>
                                    output <= "0000001110000011";
                                when others =>
                                    output <= "0000001110000011";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111000111";
                                when 1 =>
                                    output <= "0000001111000111";
                                when others =>
                                    output <= "0000001111000111";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110001011";
                                when 1 =>
                                    output <= "0000001110001011";
                                when others =>
                                    output <= "0000001110001011";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111100111";
                                when 1 =>
                                    output <= "0000001111100111";
                                when others =>
                                    output <= "0000001111100111";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001000001010";
                                when 1 =>
                                    output <= "0000001000001010";
                                when others =>
                                    output <= "0000001000001010";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000110000";
                                when 1 =>
                                    output <= "0000000000110000";
                                when others =>
                                    output <= "0000000000110000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 15 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001111100";
                                when 1 =>
                                    output <= "0000000001111100";
                                when others =>
                                    output <= "0000000001111100";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111000111";
                                when 1 =>
                                    output <= "0000001111000111";
                                when others =>
                                    output <= "0000001111000111";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001000010110";
                                when 1 =>
                                    output <= "0000001000010110";
                                when others =>
                                    output <= "0000001000010110";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001100000";
                                when 1 =>
                                    output <= "0000000001100000";
                                when others =>
                                    output <= "0000000001100000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001100010111";
                                when 1 =>
                                    output <= "0000001100010111";
                                when others =>
                                    output <= "0000001100010111";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111111011";
                                when 1 =>
                                    output <= "0000001111111011";
                                when others =>
                                    output <= "0000001111111011";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000010000000000";
                                when 1 =>
                                    output <= "0000010000000000";
                                when others =>
                                    output <= "0000010000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001011110110";
                                when 1 =>
                                    output <= "0000001011110110";
                                when others =>
                                    output <= "0000001011110110";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000011010100";
                                when 1 =>
                                    output <= "0000000011010100";
                                when others =>
                                    output <= "0000000011010100";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 16 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001001000010";
                                when 1 =>
                                    output <= "0000001001000010";
                                when others =>
                                    output <= "0000001001000010";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001100110011";
                                when 1 =>
                                    output <= "0000001100110011";
                                when others =>
                                    output <= "0000001100110011";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001000000";
                                when 1 =>
                                    output <= "0000000001000000";
                                when others =>
                                    output <= "0000000001000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000101101001";
                                when 1 =>
                                    output <= "0000000101101001";
                                when others =>
                                    output <= "0000000101101001";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110100111";
                                when 1 =>
                                    output <= "0000001110100111";
                                when others =>
                                    output <= "0000001110100111";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101101011";
                                when 1 =>
                                    output <= "0000001101101011";
                                when others =>
                                    output <= "0000001101101011";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110111101";
                                when 1 =>
                                    output <= "0000000110111101";
                                when others =>
                                    output <= "0000000110111101";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000100000";
                                when 1 =>
                                    output <= "0000000000100000";
                                when others =>
                                    output <= "0000000000100000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 17 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111101011";
                                when 1 =>
                                    output <= "0000001111101011";
                                when others =>
                                    output <= "0000001111101011";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000110000101";
                                when 1 =>
                                    output <= "0000000110000101";
                                when others =>
                                    output <= "0000000110000101";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001111100";
                                when 1 =>
                                    output <= "0000000001111100";
                                when others =>
                                    output <= "0000000001111100";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001100001111";
                                when 1 =>
                                    output <= "0000001100001111";
                                when others =>
                                    output <= "0000001100001111";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111101111";
                                when 1 =>
                                    output <= "0000001111101111";
                                when others =>
                                    output <= "0000001111101111";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001001010110";
                                when 1 =>
                                    output <= "0000001001010110";
                                when others =>
                                    output <= "0000001001010110";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000111100";
                                when 1 =>
                                    output <= "0000000000111100";
                                when others =>
                                    output <= "0000000000111100";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 18 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111111011";
                                when 1 =>
                                    output <= "0000001111111011";
                                when others =>
                                    output <= "0000001111111011";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000111111001";
                                when 1 =>
                                    output <= "0000000111111001";
                                when others =>
                                    output <= "0000000111111001";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000011001000";
                                when 1 =>
                                    output <= "0000000011001000";
                                when others =>
                                    output <= "0000000011001000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000111100001";
                                when 1 =>
                                    output <= "0000000111100001";
                                when others =>
                                    output <= "0000000111100001";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001101110011";
                                when 1 =>
                                    output <= "0000001101110011";
                                when others =>
                                    output <= "0000001101110011";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111111011";
                                when 1 =>
                                    output <= "0000001111111011";
                                when others =>
                                    output <= "0000001111111011";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111001011";
                                when 1 =>
                                    output <= "0000001111001011";
                                when others =>
                                    output <= "0000001111001011";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001000010110";
                                when 1 =>
                                    output <= "0000001000010110";
                                when others =>
                                    output <= "0000001000010110";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000111000";
                                when 1 =>
                                    output <= "0000000000111000";
                                when others =>
                                    output <= "0000000000111000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 19 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001010011010";
                                when 1 =>
                                    output <= "0000001010011010";
                                when others =>
                                    output <= "0000001010011010";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001111110111";
                                when 1 =>
                                    output <= "0000001111110111";
                                when others =>
                                    output <= "0000001111110111";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110011111";
                                when 1 =>
                                    output <= "0000001110011111";
                                when others =>
                                    output <= "0000001110011111";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001110011111";
                                when 1 =>
                                    output <= "0000001110011111";
                                when others =>
                                    output <= "0000001110011111";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000001000101110";
                                when 1 =>
                                    output <= "0000001000101110";
                                when others =>
                                    output <= "0000001000101110";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001011100";
                                when 1 =>
                                    output <= "0000000001011100";
                                when others =>
                                    output <= "0000000001011100";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 20 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000010100000";
                                when 1 =>
                                    output <= "0000000010100000";
                                when others =>
                                    output <= "0000000010100000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000001101100";
                                when 1 =>
                                    output <= "0000000001101100";
                                when others =>
                                    output <= "0000000001101100";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 21 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 22 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 23 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 24 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 25 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when 26 =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
                when others =>
                    case addressY is
                        when 0 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 1 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 2 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 3 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 4 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 5 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 6 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 7 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 8 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 9 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 10 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 11 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 12 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 13 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 14 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 15 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 16 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 17 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 18 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 19 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 20 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 21 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 22 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 23 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 24 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 25 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when 26 =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                        when others =>
                            case addressZ is
                                when 0 =>
                                    output <= "0000000000000000";
                                when 1 =>
                                    output <= "0000000000000000";
                                when others =>
                                    output <= "0000000000000000";
                            end case;
                    end case;
            end case;

        end if;
    end process;
end architecture;
